-- HOE1
