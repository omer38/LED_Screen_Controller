-- OUTPUTS HLATCH AND DATA IN SYNCHRONIZATION
