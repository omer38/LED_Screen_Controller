-- 12.5 MHZ clock
